`ifndef PRJ_DEFINES
`define PRJ_DEFINES

//`define DEBUG_HW

`define XILINX
//`define SIMULATION
//`define SPARTAN7

`define USART_EN
//`define I2C_EN
//`define HDMI_EN
//`define DDR_EN
//`define PG_EN
//`define DSI_EN
//`define PIX_READER_EN
//`define SYS_TIMER_EN

`endif