`ifndef PRJ_DEFINES
`define PRJ_DEFINES

//`define SIMULATION
`define XILINX
//`define SPARTAN7


`endif