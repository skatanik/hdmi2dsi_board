`ifndef PRJ_DEFINES
`define PRJ_DEFINES

`define XILINX
//`define SIMULATION
//`define SPARTAN7


`endif